library verilog;
use verilog.vl_types.all;
entity testebench_c is
end testebench_c;
