module testbench();

	reg [3:0]A, B;
	wire [4:0]S;

	
	somador_4bits dut (A, B, S);
	
	initial
		begin
					A = 3'b000; B = 3'b000; #50
					A = 3'b001; B = 3'b000; #50
					A = 3'b010; B = 3'b000; #50
					A = 3'b011; B = 3'b000; #50
					A = 3'b100; B = 3'b000; #50
					A = 3'b101; B = 3'b000; #50
					A = 3'b111; B = 3'b000; #50
					
					B = 3'b000; A = 3'b000; #50
					B = 3'b001; A = 3'b000; #50
					B = 3'b010; A = 3'b000; #50
					B = 3'b011; A = 3'b000; #50
					B = 3'b100; A = 3'b000; #50
					B = 3'b101; A = 3'b000; #50
					B = 3'b111; A = 3'b000; #50;
					
					A = 3'b000; B = 3'b011; #50
					A = 3'b001; B = 3'b100; #50
					A = 3'b010; B = 3'b101; #50
					B = 3'b011; A = 3'b111; #50
					B = 3'b100; A = 3'b001; #50
					B = 3'b101; A = 3'b010; #50
					B = 3'b111; A = 3'b101; #50;
			end
endmodule
