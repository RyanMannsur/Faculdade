library verilog;
use verilog.vl_types.all;
entity testebench_decodificador is
end testebench_decodificador;
